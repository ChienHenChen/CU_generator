//This delay chians element is designed for Beta version MemGen
//Version: V0
//Date: Jun 2020
//Author: Chien-Hen Chen

//-------------------------------
// Parameter definition
//-------------------------------

//-------------------------------
// Input and output definition
//-------------------------------
module DLY_MODULE (
	//Input port
	input in,
	//Output port
);

//Wire Definition
assign in0=in;

//Delay cells instantiation

//Output assign
endmodule
